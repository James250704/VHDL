library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity Final_01 is
    port (
        SW   : in STD_LOGIC_VECTOR(9 downto 0);
        LEDG : out STD_LOGIC_VECTOR(9 downto 0)
    );
end entity;

architecture Behavioral of Final_01 is
begin

end architecture;
